`timescale 1ns / 1ps

`include "../src/modules/alu.v"

module ALU_tb;

    reg [31:0] srcA;
    reg [31:0] srcB;
    reg [2:0] ALUControl;
    wire [31:0] result;

    // Instanciar la ALU
    ALU uut (
        .srcA(srcA),
        .srcB(srcB),
        .ALUControl(ALUControl),
        .result(result)
    );

    initial begin
        // Prueba de suma
        srcA = 32'd10;
        srcB = 32'd5;
        ALUControl = 3'b000; // Suma
        #10;
        
        // Prueba de resta
        ALUControl = 3'b001; // Resta
        #10;
        
        // Prueba de AND
        ALUControl = 3'b010; // AND
        #10;
        
        // Prueba de OR
        ALUControl = 3'b011; // OR
        #10;
        
        // Prueba de SLT (Set Less Than)
        srcA = 32'd5;
        srcB = 32'd10;
        ALUControl = 3'b101; // SLT
        #10;

        // Fin de la simulación
        $finish;
    end

endmodule
